package comb_gp_pkg;
  `include "comb_circuit.sv"
  `inlcude "fitness_func.sv"
endpackage