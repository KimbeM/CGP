package comb_gp_pkg;
  `include "comb_circuit.sv"
endpackage